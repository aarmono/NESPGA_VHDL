
PACKAGE ALT_CUSP_PACKAGE IS

END ALT_CUSP_PACKAGE;
